module music_player (
// TODO: fill in your implementation from lab 4!

);



endmodule